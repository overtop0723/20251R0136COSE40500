// OR Gate

module or2(x, y, o);

input x, y;
output o;

assign o=x|y;

endmodule